package scoreboard_pkg;

endpackage
