library verilog;
use verilog.vl_types.all;
entity scoreboard_pkg is
end scoreboard_pkg;
