package svm_component_pkg;
class svm_component;
endclass // svm_component_pkg
endpackage
