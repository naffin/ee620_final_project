module top;
	import lc3_interface_pkg::*;
	lc3_if lc3if
   test tb();
endmodule
