package Scoreboard_pkg;
   import Transaction_pkg::*;
class Scoreboard;
   function void compare_expected(Transaction t);
      // fill in
   endfunction
endclass

endpackage
